module m2Filler(
	input reset,
	input clk,
	input bufGetWord,
	input [7:0]bufRdPointer,
	output reg [11:0]dataWord
);

reg once2, once1;
reg [7:0]dat1012, dat6012;
always@(negedge reset or posedge clk)begin
	if (~reset) begin
		dataWord <= 0;
		dat1012 <= 0;
		dat6012 <= 0;
		once1 <= 0;
		once2 <= 0;
		dataWord <= 0;
	end else begin
		
			if(bufGetWord) begin

				case((bufRdPointer))
					0,4,8,12,16,20,24,28,32,36,40,44,48,52,56,60,64,68,72,76,80,84,88,92,96,100,104,108,112,116,120,124,128,132,136,140,144,148,152,156,160,164,168,172,176,180,184,188,192,196,200,204,208,212,216,220,224,228,232,236,240,244,248,252:
					begin // up count a10-b12
						dataWord <= {1'b0, dat1012[7:0],3'b0};
						if ((bufRdPointer == 0) || (bufRdPointer == 128)) begin
							if(once1==0)begin
								dat1012 <= dat1012 + 1'b1;
								once1=1;
							end
						end
					end
					1,5,9,13,17,21,25,29,33,37,41,45,49,53,57,61,65,69,73,77,81,85,89,93,97,101,105,109,113,117,121,125,129,133,137,141,145,149,153,157,161,165,169,173,177,181,185,189,193,197,201,205,209,213,217,221,225,229,233,237,241,245,249,253:
					begin	// down count a20-b12
						dataWord <= {1'b0, dat6012[7:0],3'b0};
						if(once2==0)begin
							dat6012 <= dat6012 - 1'b1;
							once2=1;
						end
					end
					2,6,10,14,18,22,26,30,34,38,42,46,50,54,58,62,66,70,74,78,82,86,90,94,98,102,106,110,114,118,122,126,130,134,138,142,146,150,154,158,162,166,170,174,178,182,186,190,194,198,202,206,210,214,218,222,226,230,234,238,242,246,250,254:
					begin
						dataWord <= {1'b0, 8'd111, 3'b0};
						once1=0;
						once2=0;
					end
					3,7,11,15,19,23,27,31,35,39,43,47,51,55,59,63,67,71,75,79,83,87,91,95,99,103,107,111,115,119,123,127,131,135,139,143,147,151,155,159,163,167,171,175,179,183,187,191,195,199,203,207,211,215,219,223,227,231,235,239,243,247,251,255:
					begin
						dataWord <= {1'b0, 8'd222, 3'b0};
					end
					default: dataWord <= {1'b0, 8'd0, 3'b010};
				endcase
			end

	end
end
endmodule
