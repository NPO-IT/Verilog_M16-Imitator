module m4Filler(
	input reset,
	input clk,
	input bufGetWord,
	input [8:0]bufRdPointer,
	output reg [11:0]dataWord
);

reg once2, once1;
reg [7:0]dat1012, dat6012;
always@(negedge reset or posedge clk)begin
	if (~reset) begin
		dataWord <= 0;
		dat1012 <= 0;
		dat6012 <= 0;
		once1 <= 0;
		once2 <= 0;
		dataWord <= 0;
	end else begin
		
			if(bufGetWord) begin

				case((bufRdPointer))
					0,8,16,24,32,40,48,56,64,72,80,88,96,104,112,120,128,136,144,152,160,168,176,184,192,200,208,216,224,232,240,248,256,264,272,280,288,296,304,312,320,328,336,344,352,360,368,376,384,392,400,408,416,424,432,440,448,456,464,472,480,488,496,504:
					begin // up count a10-b12
						dataWord <= {1'b0, dat1012[7:0],3'b000};
						if ((bufRdPointer == 0) || (bufRdPointer == 256)) begin
							if(once1==0)begin
								dat1012 <= dat1012 + 1'b1;
								once1=1;
							end
						end
					end
					5,13,21,29,37,45,53,61,69,77,85,93,101,109,117,125,133,141,149,157,165,173,181,189,197,205,213,221,229,237,245,253,261,269,277,285,293,301,309,317,325,333,341,349,357,365,373,381,389,397,405,413,421,429,437,445,453,461,469,477,485,493,501,509:
					begin	// down count a60-b12
						dataWord <= {1'b0, dat6012[7:0],3'b001};
						if(once2==0)begin
							dat6012 <= dat6012 - 1'b1;
							once2=1;
						end
					end
					1,9,17,25,33,41,49,57,65,73,81,89,97,105,113,121,129,137,145,153,161,169,177,185,193,201,209,217,225,233,241,249,257,265,273,281,289,297,305,313,321,329,337,345,353,361,369,377,385,393,401,409,417,425,433,441,449,457,465,473,481,489,497,505:
					begin
						dataWord <= {1'b0, 8'd11, 3'b001};
						once1=0;
					end
					2,10,18,26,34,42,50,58,66,74,82,90,98,106,114,122,130,138,146,154,162,170,178,186,194,202,210,218,226,234,242,250,258,266,274,282,290,298,306,314,322,330,338,346,354,362,370,378,386,394,402,410,418,426,434,442,450,458,466,474,482,490,498,506:
					begin
						dataWord <= {1'b0, 8'd22, 3'b000};
					end
					3,11,19,27,35,43,51,59,67,75,83,91,99,107,115,123,131,139,147,155,163,171,179,187,195,203,211,219,227,235,243,251,259,267,275,283,291,299,307,315,323,331,339,347,355,363,371,379,387,395,403,411,419,427,435,443,451,459,467,475,483,491,499,507:
					begin
						dataWord <= {1'b0, 8'd33, 3'b001};
					end
					4,12,20,28,36,44,52,60,68,76,84,92,100,108,116,124,132,140,148,156,164,172,180,188,196,204,212,220,228,236,244,252,260,268,276,284,292,300,308,316,324,332,340,348,356,364,372,380,388,396,404,412,420,428,436,444,452,460,468,476,484,492,500,508:
					begin
						dataWord <= {1'b0, 8'd44, 3'b000};
					end
					6,14,22,30,38,46,54,62,70,78,86,94,102,110,118,126,134,142,150,158,166,174,182,190,198,206,214,222,230,238,246,254,262,270,278,286,294,302,310,318,326,334,342,350,358,366,374,382,390,398,406,414,422,430,438,446,454,462,470,478,486,494,502,510:
					begin
						dataWord <= {1'b0, 8'd66, 3'b000};
						once2=0;
					end
					7,15,23,31,39,47,55,63,71,79,87,95,103,111,119,127,135,143,151,159,167,175,183,191,199,207,215,223,231,239,247,255,263,271,279,287,295,303,311,319,327,335,343,351,359,367,375,383,391,399,407,415,423,431,439,447,455,463,471,479,487,495,503,511:
					begin
						dataWord <= {1'b0, 8'd77, 3'b001};
					end
					default: dataWord <= {1'b0, 8'd0, 3'b010};
				endcase
			end

	end
end
endmodule
